library verilog;
use verilog.vl_types.all;
entity rowbuffer_vlg_vec_tst is
end rowbuffer_vlg_vec_tst;
